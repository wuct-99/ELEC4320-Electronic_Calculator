`ifndef TOP_ENV_DEF__SV
`define TOP_ENV_DEF__SV

//`define IMEM harness.u_sisyphus_core.u_sisyphus_ifu.u_imem

//parameter OPCODE_LUI    = 7'b011_0111;

`endif
