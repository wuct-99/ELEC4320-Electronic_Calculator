`ifndef CHK_INTERFACE__SV
`define CHK_INTERFACE__SV

interface chk_interface(input clk);
    //bit wrb_vld;
    //bit mem_vld;
    //bit [31:0] ireg [32];
    //bit [31:0] dmem [4][256];
    //bit [31:0] pc;
endinterface 
`endif
