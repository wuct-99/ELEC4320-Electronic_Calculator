`ifndef TC_PACKAGE__SV
`define TC_PACKAGE__SV

import uvm_pkg::*;
import cfg_package::*;
import top_env_package::*;

`endif

