module cal_top(
	//input
	clk,
	rst_n,
);

//Core input
input clk;
input rst_n;


endmodule
